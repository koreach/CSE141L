//Refer to LECTURE 7
module top(
	input clk,
		  reset,
	output logic done
	);

//You need a program counter

//InstructionROM lookup and how wide is its output. So the lookup table.

//Register file

//ALU