/*********************************************
 *  Brianna Yamanaka                         *   
 *  Jeffrey Trang                            *   
 *  Goo Gu                                   *   
 *  Byunggwan Lim                            *   
 *                                           *   
 *  CSE141L Lab3                             *   
 *                                           *   
 *  Fetch unit comprises program counter     *   
 *  and instruction memory			         *
 *                                           *   
 *********************************************/
