//do we need an instROM?


